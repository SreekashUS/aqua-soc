`include "../../regFile/regFile2R1W.v"
`include "../../branch/simple/simpleBranch.v"
`include "../../arb/tdmArbiter/tdmArbiter.v"
`include "../../core/RV32I/rv32iDecoder.v"
`include "../../core/alu/aluRv32i.v"
`include "../../"

module aqua_pygmy
#(

)
(

);

	//Default pipeline stages
	/*
	|- Fetch
	|- Decode
	|- Execute
	|- Writeback
	|- Memory access
	*/

endmodule